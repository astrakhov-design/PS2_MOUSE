//character mode LCD bitmap
//Author: Aleksander Strakhov
//Date: 05.04.2020

module LCD_character_bitmap(
	input clk,
	input [9:0] addr,
	output reg [7:0] data
	);
	
	reg [9:0] addr_reg;
	
	always @ (posedge clk)
		begin
			addr_reg <= addr;
		end
		
	always @*
		begin
			case (addr_reg)
			//code blank
			10'h000: data = 8'b0000_0000;
			10'h001: data = 8'b0000_0000;
			10'h002: data = 8'b0000_0000;
			10'h003: data = 8'b0000_0000;
			10'h004: data = 8'b0000_0000;
			10'h005: data = 8'b0000_0000;
			10'h006: data = 8'b0000_0000;
			10'h007: data = 8'b0000_0000;
			//code !
			10'h008: data = 8'b0001_1000;
			10'h009: data = 8'b0001_1000;
			10'h00a: data = 8'b0001_1000;
			10'h00b: data = 8'b0001_1000;
			10'h00c: data = 8'b0000_0000;
			10'h00d: data = 8'b0000_0000;
			10'h00e: data = 8'b0001_1000;
			10'h00f: data = 8'b0000_0000;
			//code "
			10'h010: data = 8'b0110_0110;
			10'h011: data = 8'b0110_0110;
			10'h012: data = 8'b0110_0110;
			10'h013: data = 8'b0000_0000;
			10'h014: data = 8'b0000_0000;
			10'h015: data = 8'b0000_0000;
			10'h016: data = 8'b0000_0000;
			10'h017: data = 8'b0000_0000;
			//code #
			10'h018: data = 8'b0010_0100;
			10'h019: data = 8'b0010_0100;
			10'h01a: data = 8'b1111_1111;
			10'h01b: data = 8'b0010_0100;
			10'h01c: data = 8'b1111_1111;
			10'h01d: data = 8'b0010_0100;
			10'h01e: data = 8'b0010_0100;
			10'h01f: data = 8'b0000_0000;
			//code $
			10'h020: data = 8'b0001_1000;
			10'h021: data = 8'b0011_1111;
			10'h022: data = 8'b1100_0000;
			10'h023: data = 8'b0011_1100;
			10'h024: data = 8'b0001_1011;
			10'h025: data = 8'b1111_1100;
			10'h026: data = 8'b0001_1000;
			10'h027: data = 8'b0000_0000;
			//code %
			10'h028: data = 8'b0000_0000;
			10'h029: data = 8'b0110_0010;
			10'h02a: data = 8'b0110_0100;
			10'h02b: data = 8'b0000_1000;
			10'h02c: data = 8'b0001_0000;
			10'h02d: data = 8'b0010_0110;
			10'h02e: data = 8'b0100_0110;
			10'h02f: data = 8'b0000_0000;
			//code &
			10'h030: data = 8'b0011_0000;
			10'h031: data = 8'b0100_1000;
			10'h032: data = 8'b0011_0000;
			10'h033: data = 8'b0101_0110;
			10'h034: data = 8'b1000_1000;
			10'h035: data = 8'b1000_1000;
			10'h036: data = 8'b0111_0110;
			10'h037: data = 8'b0000_0000;
			//code '
			10'h038: data = 8'b0001_0000;
			10'h039: data = 8'b0001_0000;
			10'h03a: data = 8'b0010_0000;
			10'h03b: data = 8'b0000_0000;
			10'h03c: data = 8'b0000_0000;
			10'h03d: data = 8'b0000_0000;
			10'h03e: data = 8'b0000_0000;
			10'h03f: data = 8'b0000_0000;
			//code (
			10'h040: data = 8'b0001_0000;
			10'h041: data = 8'b0010_0000;
			10'h042: data = 8'b0100_0000;
			10'h043: data = 8'b0100_0000;
			10'h044: data = 8'b0100_0000;
			10'h045: data = 8'b0010_0000;
			10'h046: data = 8'b0001_0000;
			10'h047: data = 8'b0000_0000;
			//code )
			10'h048: data = 8'b0010_0000;
			10'h049: data = 8'b0001_0000;
			10'h04a: data = 8'b0000_1000;
			10'h04b: data = 8'b0000_1000;
			10'h04c: data = 8'b0000_1000;
			10'h04d: data = 8'b0001_0000;
			10'h04e: data = 8'b0010_0000;
			10'h04f: data = 8'b0000_0000;
			//code *
			10'h050: data = 8'b0000_0000;
			10'h051: data = 8'b0100_0100;
			10'h052: data = 8'b0011_1000;
			10'h053: data = 8'b1111_1110;
			10'h054: data = 8'b0011_1000;
			10'h055: data = 8'b0100_0100;
			10'h056: data = 8'b0000_0000;
			10'h057: data = 8'b0000_0000;
			// code +
			10'h058: data = 8'b0000_0000;
			10'h059: data = 8'b0001_0000;
			10'h05a: data = 8'b0001_0000;
			10'h05b: data = 8'b0111_1100;
			10'h05c: data = 8'b0001_0000;
			10'h05d: data = 8'b0001_0000;
			10'h05e: data = 8'b0000_0000;
			10'h05f: data = 8'b0000_0000;
			// code ,
			10'h060: data = 8'b0000_0000;
			10'h061: data = 8'b0000_0000;
			10'h062: data = 8'b0000_0000;
			10'h063: data = 8'b0000_0000;
			10'h064: data = 8'b0001_0000;
			10'h065: data = 8'b0001_0000;
			10'h066: data = 8'b0010_0000;
			10'h067: data = 8'b0000_0000;
			// code -
			10'h068: data = 8'b0000_0000;
			10'h069: data = 8'b0000_0000;
			10'h06a: data = 8'b0000_0000;
			10'h06b: data = 8'b0111_1110;
			10'h06c: data = 8'b0000_0000;
			10'h06d: data = 8'b0000_0000;
			10'h06e: data = 8'b0000_0000;
			10'h06f: data = 8'b0000_0000;
			// code .
			10'h070: data = 8'b0000_0000;
			10'h071: data = 8'b0000_0000;
			10'h072: data = 8'b0000_0000;
			10'h073: data = 8'b0000_0000;
			10'h074: data = 8'b0000_0000;
			10'h075: data = 8'b0001_0000;
			10'h076: data = 8'b0001_0000;
			10'h077: data = 8'b0000_0000;
			// code /
			10'h078: data = 8'b0000_0000;
			10'h079: data = 8'b0000_0010;
			10'h07a: data = 8'b0000_0100;
			10'h07b: data = 8'b0000_1000;
			10'h07c: data = 8'b0001_0000;
			10'h07d: data = 8'b0010_0000;
			10'h07e: data = 8'b0100_0000;
			10'h07f: data = 8'b0000_0000;
			// code 0
			10'h080: data = 8'b0111_1100;
			10'h081: data = 8'b1100_0110;
			10'h082: data = 8'b1100_0110;
			10'h083: data = 8'b1101_0110;
			10'h084: data = 8'b1100_0110;
			10'h085: data = 8'b1100_0110;
			10'h086: data = 8'b0111_1100;
			10'h087: data = 8'b0000_0000;
			// code 1
			10'h088: data = 8'b0011_0000;
			10'h089: data = 8'b0111_0000;
			10'h08a: data = 8'b0011_0000;
			10'h08b: data = 8'b0011_0000;
			10'h08c: data = 8'b0011_0000;
			10'h08d: data = 8'b0011_0000;
			10'h08e: data = 8'b1111_1100;
			10'h08f: data = 8'b0000_0000;
			//code 2
			10'h090: data = 8'b0111_1000;
			10'h091: data = 8'b1100_1100;
			10'h092: data = 8'b0000_1100;
			10'h093: data = 8'b0011_1000;
			10'h094: data = 8'b0110_0000;
			10'h095: data = 8'b1100_0011;
			10'h096: data = 8'b1111_1100;
			10'h097: data = 8'b0000_0000;
			// code 3
			10'h098: data = 8'b0111_1000;
			10'h099: data = 8'b1100_1100;
			10'h09a: data = 8'b0000_1100;
			10'h09b: data = 8'b0011_1000;
			10'h09c: data = 8'b0000_1100;
			10'h09d: data = 8'b1100_1100;
			10'h09e: data = 8'b0111_1000;
			10'h09f: data = 8'b0000_0000;
			// code 4
			10'h0a0: data = 8'b0000_0110;
			10'h0a1: data = 8'b0000_1110;
			10'h0a2: data = 8'b0001_1110;
			10'h0a3: data = 8'b0110_0110;
			10'h0a4: data = 8'b0111_1111;
			10'h0a5: data = 8'b0000_0110;
			10'h0a6: data = 8'b0000_0110;
			10'h0a7: data = 8'b0000_0000;
			// code 5
			10'h0a8: data = 8'b0111_1110;
			10'h0a9: data = 8'b0110_0000;
			10'h0aa: data = 8'b0111_1100;
			10'h0ab: data = 8'b0000_0110;
			10'h0ac: data = 8'b0000_0110;
			10'h0ad: data = 8'b0110_0110;
			10'h0ae: data = 8'b0011_1100;
			10'h0af: data = 8'b0000_0000;
			// code 6
			10'h0b0: data = 8'b0011_1100;
			10'h0b1: data = 8'b0110_0110;
			10'h0b2: data = 8'b0110_0000;
			10'h0b3: data = 8'b0111_1100;
			10'h0b4: data = 8'b0110_0110;
			10'h0b5: data = 8'b0110_0110;
			10'h0b6: data = 8'b0011_1100;
			10'h0b7: data = 8'b0000_0000;
			// code 7
			10'h0b8: data = 8'b0111_1110;
			10'h0b9: data = 8'b0110_0110;
			10'h0ba: data = 8'b0000_1100;
			10'h0bb: data = 8'b0001_1000;
			10'h0bc: data = 8'b0001_1000;
			10'h0bd: data = 8'b0001_1000;
			10'h0be: data = 8'b0001_1000;
			10'h0bf: data = 8'b0000_0000;
			// code 8
			10'h0c0: data = 8'b0011_1100;
			10'h0c1: data = 8'b0110_0110;
			10'h0c2: data = 8'b0110_0110;
			10'h0c3: data = 8'b0011_1100;
			10'h0c4: data = 8'b0110_0110;
			10'h0c5: data = 8'b0110_0110;
			10'h0c6: data = 8'b0011_1100;
			10'h0c7: data = 8'b0000_0000;
			// code 9
			10'h0c8: data = 8'b0011_1100;
			10'h0c9: data = 8'b0110_0110;
			10'h0ca: data = 8'b0110_0110;
			10'h0cb: data = 8'b0011_1110;
			10'h0cc: data = 8'b0000_0110;
			10'h0cd: data = 8'b0110_0110;
			10'h0ce: data = 8'b0011_1100;
			10'h0cf: data = 8'b0000_0000;
			//code :
			10'h0d0: data = 8'b0000_0000;
			10'h0d1: data = 8'b0000_0000;
			10'h0d2: data = 8'b0001_1000;
			10'h0d3: data = 8'b0000_0000;
			10'h0d4: data = 8'b0000_0000;
			10'h0d5: data = 8'b0001_1000;
			10'h0d6: data = 8'b0000_0000;
			10'h0d7: data = 8'b0000_0000;
			//code ;
			10'h0d8: data = 8'b0000_0000;
			10'h0d9: data = 8'b0000_0000;
			10'h0da: data = 8'b0001_1000;
			10'h0db: data = 8'b0000_0000;
			10'h0dc: data = 8'b0000_0000;
			10'h0dd: data = 8'b0001_1000;
			10'h0de: data = 8'b0001_1000;
			10'h0df: data = 8'b0011_0000;
			// code <
			10'h0e0: data = 8'b0000_1110;
			10'h0e1: data = 8'b0001_1000;
			10'h0e2: data = 8'b0011_0000;
			10'h0e3: data = 8'b0110_0000;
			10'h0e4: data = 8'b0011_0000;
			10'h0e5: data = 8'b0001_1000;
			10'h0e6: data = 8'b0000_1110;
			10'h0e7: data = 8'b0000_0000;
			// code =
			10'h0e8: data = 8'b0000_0000;
			10'h0e9: data = 8'b0000_0000;
			10'h0ea: data = 8'b0111_1110;
			10'h0eb: data = 8'b0000_0000;
			10'h0ec: data = 8'b0111_1110;
			10'h0ed: data = 8'b0000_0000;
			10'h0ee: data = 8'b0000_0000;
			10'h0ef: data = 8'b0000_0000;
			//code >
			10'h0f0: data = 8'b0111_0000;
			10'h0f1: data = 8'b0001_1000;
			10'h0f2: data = 8'b0000_1100;
			10'h0f3: data = 8'b0000_0110;
			10'h0f4: data = 8'b0000_1100;
			10'h0f5: data = 8'b0001_1000;
			10'h0f6: data = 8'b0111_0000;
			10'h0f7: data = 8'b0000_0000;
			// code ?
			10'h0f8: data = 8'b0011_1100;
			10'h0f9: data = 8'b0110_0110;
			10'h0fa: data = 8'b0000_0110;
			10'h0fb: data = 8'b0000_1100;
			10'h0fc: data = 8'b0001_1000;
			10'h0fd: data = 8'b0000_0000;
			10'h0fe: data = 8'b0001_1000;
			10'h0ff: data = 8'b0000_0000;
			//code @
			10'h100: data = 8'b0011_1100;
			10'h101: data = 8'b0110_0110;
			10'h102: data = 8'b0110_1110;
			10'h103: data = 8'b0110_1110;
			10'h104: data = 8'b0110_0000;
			10'h105: data = 8'b0110_0110;
			10'h106: data = 8'b0011_1100;
			10'h107: data = 8'b0000_0000;
			//code A
			10'h108: data = 8'b0001_1000;
			10'h109: data = 8'b0011_1100;
			10'h10a: data = 8'b0110_0110;
			10'h10b: data = 8'b0111_1110;
			10'h10c: data = 8'b0110_0110;
			10'h10d: data = 8'b0110_0110;
			10'h10e: data = 8'b0110_0110;
			10'h10f: data = 8'b0000_0000;
			// code B
			10'h110: data = 8'b0111_1100;
			10'h111: data = 8'b0110_0110;
			10'h112: data = 8'b0110_0110;
			10'h113: data = 8'b0111_1100;
			10'h114: data = 8'b0110_0110;
			10'h115: data = 8'b0110_0110;
			10'h116: data = 8'b0111_1100;
			10'h117: data = 8'b0000_0000;
			//code C
			10'h118: data = 8'b0011_1100;
			10'h119: data = 8'b0110_0110;
			10'h11a: data = 8'b0110_0000;
			10'h11b: data = 8'b0110_0000;
			10'h11c: data = 8'b0110_0000;
			10'h11d: data = 8'b0110_0110;
			10'h11e: data = 8'b0011_1100;
			10'h11f: data = 8'b0000_0000;
			//code D
			10'h120: data = 8'b0111_1000;
			10'h121: data = 8'b0110_1100;
			10'h122: data = 8'b0110_0110;
			10'h123: data = 8'b0110_0110;
			10'h124: data = 8'b0110_0110;
			10'h125: data = 8'b0110_1100;
			10'h126: data = 8'b0111_1000;
			10'h127: data = 8'b0000_0000;
			//code E
			10'h128: data = 8'b0111_1110;
			10'h129: data = 8'b0110_0000;
			10'h12a: data = 8'b0110_0000;
			10'h12b: data = 8'b0111_1000;
			10'h12c: data = 8'b0110_0000;
			10'h12d: data = 8'b0110_0000;
			10'h12e: data = 8'b0111_1110;
			10'h12f: data = 8'b0000_0000;
			//code F
			10'h130: data = 8'b0111_1110;
			10'h131: data = 8'b0110_0000;
			10'h132: data = 8'b0110_0000;
			10'h133: data = 8'b0111_1000;
			10'h134: data = 8'b0110_0000;
			10'h135: data = 8'b0110_0000;
			10'h136: data = 8'b0110_0000;
			10'h137: data = 8'b0000_0000;
			//code G
			10'h138: data = 8'b0011_1100;
			10'h139: data = 8'b0110_0110;
			10'h13a: data = 8'b0110_0000;
			10'h13b: data = 8'b0110_1110;
			10'h13c: data = 8'b0110_0110;
			10'h13d: data = 8'b0110_0110;
			10'h13e: data = 8'b0011_1100;
			10'h13f: data = 8'b0000_0000;
			//code H
			10'h140: data = 8'b0110_0110;
			10'h141: data = 8'b0110_0110;
			10'h142: data = 8'b0110_0110;
			10'h143: data = 8'b0111_1110;
			10'h144: data = 8'b0110_0110;
			10'h145: data = 8'b0110_0110;
			10'h146: data = 8'b0110_0110;
			10'h147: data = 8'b0000_0000;
			//code I
			10'h148: data = 8'b0011_1100;
			10'h149: data = 8'b0001_1000;
			10'h14a: data = 8'b0001_1000;
			10'h14b: data = 8'b0001_1000;
			10'h14c: data = 8'b0001_1000;
			10'h14d: data = 8'b0001_1000;
			10'h14e: data = 8'b0011_1100;
			10'h14f: data = 8'b0000_0000;
			//code J
			10'h150: data = 8'b0001_1110;
			10'h151: data = 8'b0000_1100;
			10'h152: data = 8'b0000_1100;
			10'h153: data = 8'b0000_1100;
			10'h154: data = 8'b0000_1100;
			10'h155: data = 8'b0110_1100;
			10'h156: data = 8'b0011_1000;
			10'h157: data = 8'b0000_0000;
			//code K
			10'h158: data = 8'b0110_0110;
			10'h159: data = 8'b0110_1100;
			10'h15a: data = 8'b0111_1000;
			10'h15b: data = 8'b0111_0000;
			10'h15c: data = 8'b0111_1000;
			10'h15d: data = 8'b0110_1100;
			10'h15e: data = 8'b0110_0110;
			10'h15f: data = 8'b0000_0000;
			//code L
			10'h160: data = 8'b0110_0000;
			10'h161: data = 8'b0110_0000;
			10'h162: data = 8'b0110_0000;
			10'h163: data = 8'b0110_0000;
			10'h164: data = 8'b0110_0000;
			10'h165: data = 8'b0110_0000;
			10'h166: data = 8'b0111_1110;
			10'h167: data = 8'b0000_0000;
			//code M
			10'h168: data = 8'b0110_0011;
			10'h169: data = 8'b0111_0111;
			10'h16a: data = 8'b0111_1111;
			10'h16b: data = 8'b0110_1011;
			10'h16c: data = 8'b0110_0011;
			10'h16d: data = 8'b0110_0011;
			10'h16e: data = 8'b0110_0011;
			10'h16f: data = 8'b0000_0000;
			//code N
			10'h170: data = 8'b0110_0110;
			10'h171: data = 8'b0111_0110;
			10'h172: data = 8'b0111_1110;
			10'h173: data = 8'b0111_1110;
			10'h174: data = 8'b0110_1110;
			10'h175: data = 8'b0110_0110;
			10'h176: data = 8'b0110_0110;
			10'h177: data = 8'b0000_0000;
			//code O
			10'h178: data = 8'b0011_1100;
			10'h179: data = 8'b0110_0110;
			10'h17a: data = 8'b0110_0110;
			10'h17b: data = 8'b0110_0110;
			10'h17c: data = 8'b0110_0110;
			10'h17d: data = 8'b0110_0110;
			10'h17e: data = 8'b0011_1100;
			10'h17f: data = 8'b0000_0000;
			//code P
			10'h180: data = 8'b0111_1100;
			10'h181: data = 8'b0110_0110;
			10'h182: data = 8'b0110_0110;
			10'h183: data = 8'b0111_1100;
			10'h184: data = 8'b0110_0000;
			10'h185: data = 8'b0110_0000;
			10'h186: data = 8'b0110_0000;
			10'h187: data = 8'b0000_0000;
			//code Q
			10'h188: data = 8'b0011_1100;
			10'h189: data = 8'b0110_0110;
			10'h18a: data = 8'b0110_0110;
			10'h18b: data = 8'b0110_0110;
			10'h18c: data = 8'b0110_0110;
			10'h18d: data = 8'b0011_1100;
			10'h18e: data = 8'b0000_1110;
			10'h18f: data = 8'b0000_0000;
			//code R
			10'h190: data = 8'b0111_1100;
			10'h191: data = 8'b0110_0110;
			10'h192: data = 8'b0110_0110;
			10'h193: data = 8'b0111_1100;
			10'h194: data = 8'b0111_1000;
			10'h195: data = 8'b0110_1100;
			10'h196: data = 8'b0110_0110;
			10'h197: data = 8'b0000_0000;
			//code S
			10'h198: data = 8'b0011_1100;
			10'h199: data = 8'b0110_0110;
			10'h19a: data = 8'b0110_0000;
			10'h19b: data = 8'b0011_1100;
			10'h19c: data = 8'b0000_0110;
			10'h19d: data = 8'b0110_0110;
			10'h19e: data = 8'b0011_1100;
			10'h19f: data = 8'b0000_0000;
			//code T
			10'h1a0: data = 8'b0111_1110;
			10'h1a1: data = 8'b0001_1000;
			10'h1a2: data = 8'b0001_1000;
			10'h1a3: data = 8'b0001_1000;
			10'h1a4: data = 8'b0001_1000;
			10'h1a5: data = 8'b0001_1000;
			10'h1a6: data = 8'b0001_1000;
			10'h1a7: data = 8'b0000_0000;
			//code U
			10'h1a8: data = 8'b0110_0110;
			10'h1a9: data = 8'b0110_0110;
			10'h1aa: data = 8'b0110_0110;
			10'h1ab: data = 8'b0110_0110;
			10'h1ac: data = 8'b0110_0110;
			10'h1ad: data = 8'b0110_0110;
			10'h1ae: data = 8'b0011_1100;
			10'h1af: data = 8'b0000_0000;
			//code V
			10'h1b0: data = 8'b0110_0110;
			10'h1b1: data = 8'b0110_0110;
			10'h1b2: data = 8'b0110_0110;
			10'h1b3: data = 8'b0110_0110;
			10'h1b4: data = 8'b0110_0110;
			10'h1b5: data = 8'b0011_1100;
			10'h1b6: data = 8'b0001_1000;
			10'h1b7: data = 8'b0000_0000;
			//code W
			10'h1b8: data = 8'b0110_0011;
			10'h1b9: data = 8'b0110_0011;
			10'h1ba: data = 8'b0110_0011;
			10'h1bb: data = 8'b0110_1011;
			10'h1bc: data = 8'b0111_1111;
			10'h1bd: data = 8'b0111_0111;
			10'h1be: data = 8'b0110_0011;
			10'h1bf: data = 8'b0000_0000;
			//code X
			10'h1c0: data = 8'b0110_0110;
			10'h1c1: data = 8'b0110_0110;
			10'h1c2: data = 8'b0011_1100;
			10'h1c3: data = 8'b0001_1000;
			10'h1c4: data = 8'b0011_1100;
			10'h1c5: data = 8'b0110_0110;
			10'h1c6: data = 8'b0110_0110;
			10'h1c7: data = 8'b0000_0000;
			//code Y
			10'h1c8: data = 8'b0110_0110;
			10'h1c9: data = 8'b0110_0110;
			10'h1ca: data = 8'b0110_0110;
			10'h1cb: data = 8'b0011_1100;
			10'h1cc: data = 8'b0001_1000;
			10'h1cd: data = 8'b0001_1000;
			10'h1ce: data = 8'b0001_1000;
			10'h1cf: data = 8'b0000_0000;
			//code Z
			10'h1d0: data = 8'b0111_1110;
			10'h1d1: data = 8'b0000_0110;
			10'h1d2: data = 8'b0000_1100;
			10'h1d3: data = 8'b0001_1000;
			10'h1d4: data = 8'b0011_0000;
			10'h1d5: data = 8'b0110_0000;
			10'h1d6: data = 8'b0111_1110;
			10'h1d7: data = 8'b0000_0000;
			
			default: data = 8'b0000_0000;
			
			endcase
		end
endmodule