//character mode LCD bitmap
//Author: Aleksander Strakhov
//Date: 05.04.2020

module LCD_character_bitmap(
	input clk,
	input [9:0] addr,
	output reg [7:0] data
	);
	
	reg [9:0] addr_reg;
	
	always @ (posedge clk)
		begin
			addr_reg <= addr;
		end
		
	always @*
		begin
			case (addr_reg)
			//code blank
			10'h000: data = 8'b0000_0000;
			10'h001: data = 8'b0000_0000;
			10'h002: data = 8'b0000_0000;
			10'h003: data = 8'b0000_0000;
			10'h004: data = 8'b0000_0000;
			10'h005: data = 8'b0000_0000;
			10'h006: data = 8'b0000_0000;
			10'h007: data = 8'b0000_0000;
			//code !
			10'h008: data = 8'b0001_1000;
			10'h009: data = 8'b0001_1000;
			10'h00a: data = 8'b0001_1000;
			10'h00b: data = 8'b0001_1000;
			10'h00c: data = 8'b0000_0000;
			10'h00d: data = 8'b0000_0000;
			10'h00e: data = 8'b0001_1000;
			10'h00f: data = 8'b0000_0000;
			//code "
			10'h010: data = 8'b0110_0110;
			10'h011: data = 8'b0110_0110;
			10'h012: data = 8'b0110_0110;
			10'h013: data = 8'b0000_0000;
			10'h014: data = 8'b0000_0000;
			10'h015: data = 8'b0000_0000;
			10'h016: data = 8'b0000_0000;
			10'h017: data = 8'b0000_0000;
			//code #
			10'h018: data = 8'b0010_0100;
			10'h019: data = 8'b0010_0100;
			10'h01a: data = 8'b1111_1111;
			10'h01b: data = 8'b0010_0100;
			10'h01c: data = 8'b1111_1111;
			10'h01d: data = 8'b0010_0100;
			10'h01e: data = 8'b0010_0100;
			10'h01f: data = 8'b0000_0000;
			//code $
			10'h020: data = 8'b0001_1000;
			10'h021: data = 8'b0011_1111;
			10'h022: data = 8'b1100_0000;
			10'h023: data = 8'b0011_1100;
			10'h024: data = 8'b0001_1011;
			10'h025: data = 8'b1111_1100;
			10'h026: data = 8'b0001_1000;
			10'h027: data = 8'b0000_0000;
			//code %
			10'h028: data = 8'b0000_0000;
			10'h029: data = 8'b0110_0010;
			10'h02a: data = 8'b0110_0100;
			10'h02b: data = 8'b0000_1000;
			10'h02c: data = 8'b0001_0000;
			10'h02d: data = 8'b0010_0110;
			10'h02e: data = 8'b0100_0110;
			10'h02f: data = 8'b0000_0000;
			//code &
			10'h030: data = 8'b0011_0000;
			10'h031: data = 8'b0100_1000;
			10'h032: data = 8'b0011_0000;
			10'h033: data = 8'b0101_0110;
			10'h034: data = 8'b1000_1000;
			10'h035: data = 8'b1000_1000;
			10'h036: data = 8'b0111_0110;
			10'h037: data = 8'b0000_0000;
			//code '
			10'h038: data = 8'b0001_0000;
			10'h039: data = 8'b0001_0000;
			10'h03a: data = 8'b0010_0000;
			10'h03b: data = 8'b0000_0000;
			10'h03c: data = 8'b0000_0000;
			10'h03d: data = 8'b0000_0000;
			10'h03e: data = 8'b0000_0000;
			10'h03f: data = 8'b0000_0000;
			//code (
			10'h040: data = 8'b0001_0000;
			10'h041: data = 8'b0010_0000;
			10'h042: data = 8'b0100_0000;
			10'h043: data = 8'b0100_0000;
			10'h044: data = 8'b0100_0000;
			10'h045: data = 8'b0010_0000;
			10'h046: data = 8'b0001_0000;
			10'h047: data = 8'b0000_0000;
			//code )
			10'h048: data = 8'b0010_0000;
			10'h049: data = 8'b0001_0000;
			10'h04a: data = 8'b0000_1000;
			10'h04b: data = 8'b0000_1000;
			10'h04c: data = 8'b0000_1000;
			10'h04d: data = 8'b0001_0000;
			10'h04e: data = 8'b0010_0000;
			10'h04f: data = 8'b0000_0000;
			//code *
			10'h050: data = 8'b0000_0000;
			10'h051: data = 8'b0100_0100;
			10'h052: data = 8'b0011_1000;
			10'h053: data = 8'b1111_1110;
			10'h054: data = 8'b0011_1000;
			10'b055: data = 8'b0100_0100;
			10'b056: data = 8'b0000_0000;
			10'b057: data = 8'b0000_0000;
			// code +
			10'h058: data = 8'b0000_0000;
			10'h059: data = 8'b0001_0000;
			10'h05a: data = 8'b0001_0000;
			10'h05b: data = 8'b0111_1100;
			10'h05c: data = 8'b0001_0000;
			10'h05d: data = 8'b0001_0000;
			10'h05e: data = 8'b0000_0000;
			10'h05f: data = 8'b0000_0000;
			// code ,
			10'h060: data = 8'b0000_0000;
			10'h061: data = 8'b0000_0000;
			10'h062: data = 8'b0000_0000;
			10'h063: data = 8'b0000_0000;
			10'h064: data = 8'b0001_0000;
			10'h065: data = 8'b0001_0000;
			10'h066: data = 8'b0010_0000;
			10'h067: data = 8'b0000_0000;
			// code -
			10'h068: data = 8'b0000_0000;
			10'h069: data = 8'b0000_0000;
			10'h06a: data = 8'b0000_0000;
			10'h06b: data = 8'b0111_1110;
			10'h06c: data = 8'b0000_0000;
			10'h06d: data = 8'b0000_0000;
			10'h06e: data = 8'b0000_0000;
			10'h06f: data = 8'b0000_0000;
			// code .
			10'h070: data = 8'b0000_0000;
			10'h071: data = 8'b0000_0000;
			10'h072: data = 8'b0000_0000;
			10'h073: data = 8'b0000_0000;
			10'h074: data = 8'b0000_0000;
			10'h075: data = 8'b0001_0000;
			10'h076: data = 8'b0001_0000;
			10'h077: data = 8'b0000_0000;
			// code /
			10'h078: data = 8'b0000_0000;
			10'h079: data = 8'b0000_0010;
			10'h07a: data = 8'b0000_0100;
			10'h07b: data = 8'b0000_1000;
			10'h07c: data = 8'b0001_0000;
			10'h07d: data = 8'b0010_0000;
			10'h07e: data = 8'b0100_0000;
			10'h07f: data = 8'b0000_0000;
			// code 0
			10'h080: data = 8'b0111_1100;
			10'h081: data = 8'b1100_0110;
			10'h082: data = 8'b1100_0110;
			10'h083: data = 8'b1101_0110;
			10'h084: data = 8'b1100_0110;
			10'h085: data = 8'b1100_0110;
			10'h086: data = 8'b0111_1100;
			10'h087: data = 8'b0000_0000;
			// code 1
			10'h088: data = 8'b0011_0000;
			10'h089: data = 8'b0111_0000;
			10'h08a: data = 8'b0011_0000;
			10'h08b: data = 8'b0011_0000;
			10'h08c: data = 8'b0011_0000;
			10'h08d: data = 8'b0011_0000;
			10'h08e: data = 8'b1111_1100;
			10'h08f: data = 8'b0000_0000;
			//code 2
			10'h090: data = 8'b0111_1000;
			10'h091: data = 8'b1100_1100;
			10'h092: data = 8'b0000_1100;
			10'h093: data = 8'b0011_1000;
			10'h094: data = 8'b0110_0000;
			10'h095: data = 8'b1100_0011;
			10'h096: data = 8'b1111_1100;
			10'h097: data = 8'b0000_0000;
			// code 3
			10'h098: data = 8'b0111_1000;
			10'h099: data = 8'b1100_1100;
			10'h09a: data = 8'b0000_1100;
			10'h09b: data = 8'b0011_1000;
			10'h09c: data = 8'b0000_1100;
			10'h09d: data = 8'b1100_1100;
			10'h09e: data = 8'b0111_1000;
			10'h09f: data = 8'b0000_0000;